library verilog;
use verilog.vl_types.all;
entity tb_sys_level is
end tb_sys_level;
