library verilog;
use verilog.vl_types.all;
entity decoder is
    port(
        iCLOCK          : in     vl_logic;
        inRESET         : in     vl_logic;
        iFREE_DEFAULT   : in     vl_logic;
        iPREVIOUS_INST_VALID: in     vl_logic;
        iPREVIOUS_FAULT_PAGEFAULT: in     vl_logic;
        iPREVIOUS_FAULT_PRIVILEGE_ERROR: in     vl_logic;
        iPREVIOUS_FAULT_INVALID_INST: in     vl_logic;
        iPREVIOUS_PAGING_ENA: in     vl_logic;
        iPREVIOUS_KERNEL_ACCESS: in     vl_logic;
        iPREVIOUS_BRANCH_PREDICT: in     vl_logic;
        iPREVIOUS_BRANCH_PREDICT_ADDR: in     vl_logic_vector(31 downto 0);
        iPREVIOUS_INST  : in     vl_logic_vector(31 downto 0);
        iPREVIOUS_PC    : in     vl_logic_vector(31 downto 0);
        oPREVIOUS_LOCK  : out    vl_logic;
        oNEXT_VALID     : out    vl_logic;
        oNEXT_FAULT_PAGEFAULT: out    vl_logic;
        oNEXT_FAULT_PRIVILEGE_ERROR: out    vl_logic;
        oNEXT_FAULT_INVALID_INST: out    vl_logic;
        oNEXT_PAGING_ENA: out    vl_logic;
        oNEXT_KERNEL_ACCESS: out    vl_logic;
        oNEXT_BRANCH_PREDICT: out    vl_logic;
        oNEXT_BRANCH_PREDICT_ADDR: out    vl_logic_vector(31 downto 0);
        oNEXT_SOURCE0_ACTIVE: out    vl_logic;
        oNEXT_SOURCE1_ACTIVE: out    vl_logic;
        oNEXT_SOURCE0_SYSREG: out    vl_logic;
        oNEXT_SOURCE1_SYSREG: out    vl_logic;
        oNEXT_SOURCE0_SYSREG_RENAME: out    vl_logic;
        oNEXT_SOURCE1_SYSREG_RENAME: out    vl_logic;
        oNEXT_ADV_ACTIVE: out    vl_logic;
        oNEXT_DESTINATION_SYSREG: out    vl_logic;
        oNEXT_DEST_RENAME: out    vl_logic;
        oNEXT_WRITEBACK : out    vl_logic;
        oNEXT_FLAGS_WRITEBACK: out    vl_logic;
        oNEXT_FRONT_COMMIT_WAIT: out    vl_logic;
        oNEXT_CMD       : out    vl_logic_vector(4 downto 0);
        oNEXT_CC_AFE    : out    vl_logic_vector(3 downto 0);
        oNEXT_SOURCE0   : out    vl_logic_vector(4 downto 0);
        oNEXT_SOURCE1   : out    vl_logic_vector(31 downto 0);
        oNEXT_ADV_DATA  : out    vl_logic_vector(5 downto 0);
        oNEXT_SOURCE0_FLAGS: out    vl_logic;
        oNEXT_SOURCE1_IMM: out    vl_logic;
        oNEXT_DESTINATION: out    vl_logic_vector(4 downto 0);
        oNEXT_EX_SYS_REG: out    vl_logic;
        oNEXT_EX_SYS_LDST: out    vl_logic;
        oNEXT_EX_LOGIC  : out    vl_logic;
        oNEXT_EX_SHIFT  : out    vl_logic;
        oNEXT_EX_ADDER  : out    vl_logic;
        oNEXT_EX_MUL    : out    vl_logic;
        oNEXT_EX_SDIV   : out    vl_logic;
        oNEXT_EX_UDIV   : out    vl_logic;
        oNEXT_EX_LDST   : out    vl_logic;
        oNEXT_EX_BRANCH : out    vl_logic;
        oNEXT_PC        : out    vl_logic_vector(31 downto 0);
        iNEXT_LOCK      : in     vl_logic
    );
end decoder;
