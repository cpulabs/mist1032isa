library verilog;
use verilog.vl_types.all;
entity core_debug is
    port(
        iCLOCK          : in     vl_logic;
        inRESET         : in     vl_logic;
        iCMD_REQ        : in     vl_logic;
        oCMD_BUSY       : out    vl_logic;
        iCMD_COMMAND    : in     vl_logic_vector(3 downto 0);
        iCMD_TARGET     : in     vl_logic_vector(7 downto 0);
        iCMD_DATA       : in     vl_logic_vector(31 downto 0);
        oRESP_VALID     : out    vl_logic;
        oRESP_ERROR     : out    vl_logic;
        oRESP_DATA      : out    vl_logic_vector(31 downto 0);
        oDEBUG_CORE_REQ : out    vl_logic;
        oDEBUG_CORE_STOP: out    vl_logic;
        oDEBUG_CORE_START: out    vl_logic;
        iDEBUG_CORE_ACK : in     vl_logic;
        iREG_R_GR0      : in     vl_logic_vector(31 downto 0);
        iREG_R_GR1      : in     vl_logic_vector(31 downto 0);
        iREG_R_GR2      : in     vl_logic_vector(31 downto 0);
        iREG_R_GR3      : in     vl_logic_vector(31 downto 0);
        iREG_R_GR4      : in     vl_logic_vector(31 downto 0);
        iREG_R_GR5      : in     vl_logic_vector(31 downto 0);
        iREG_R_GR6      : in     vl_logic_vector(31 downto 0);
        iREG_R_GR7      : in     vl_logic_vector(31 downto 0);
        iREG_R_GR8      : in     vl_logic_vector(31 downto 0);
        iREG_R_GR9      : in     vl_logic_vector(31 downto 0);
        iREG_R_GR10     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR11     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR12     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR13     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR14     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR15     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR16     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR17     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR18     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR19     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR20     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR21     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR22     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR23     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR24     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR25     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR26     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR27     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR28     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR29     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR30     : in     vl_logic_vector(31 downto 0);
        iREG_R_GR31     : in     vl_logic_vector(31 downto 0);
        iREG_R_CPUIDR   : in     vl_logic_vector(31 downto 0);
        iREG_R_TIDR     : in     vl_logic_vector(31 downto 0);
        iREG_R_FLAGR    : in     vl_logic_vector(31 downto 0);
        iREG_R_PCR      : in     vl_logic_vector(31 downto 0);
        iREG_R_SPR      : in     vl_logic_vector(31 downto 0);
        iREG_R_PSR      : in     vl_logic_vector(31 downto 0);
        iREG_R_IOSAR    : in     vl_logic_vector(31 downto 0);
        iREG_R_TISR     : in     vl_logic_vector(31 downto 0);
        iREG_R_IDTR     : in     vl_logic_vector(31 downto 0);
        iREG_R_FI0R     : in     vl_logic_vector(31 downto 0);
        iREG_R_FI1R     : in     vl_logic_vector(31 downto 0);
        iREG_R_FRCLR    : in     vl_logic_vector(31 downto 0);
        iREG_R_FRCHR    : in     vl_logic_vector(31 downto 0);
        iREG_R_PTIDR    : in     vl_logic_vector(31 downto 0);
        iREG_R_PFLAGR   : in     vl_logic_vector(31 downto 0);
        iREG_R_PPCR     : in     vl_logic_vector(31 downto 0);
        iREG_R_PPSR     : in     vl_logic_vector(31 downto 0);
        iREG_R_PPDTR    : in     vl_logic_vector(31 downto 0)
    );
end core_debug;
