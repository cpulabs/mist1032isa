library verilog;
use verilog.vl_types.all;
entity exception_manager is
    port(
        iCLOCK          : in     vl_logic;
        inRESET         : in     vl_logic;
        oFREE_REGISTER_LOCK: out    vl_logic;
        oFREE_PIPELINE_STOP: out    vl_logic;
        oFREE_REFRESH   : out    vl_logic;
        oFREE_RESTART   : out    vl_logic;
        oFREE_PC_SET    : out    vl_logic;
        oFREE_PC        : out    vl_logic_vector(31 downto 0);
        oFREE_PPCR_SET  : out    vl_logic;
        oFREE_PPCR      : out    vl_logic_vector(31 downto 0);
        oFREE_FI0R_SET  : out    vl_logic;
        oFREE_FI0R      : out    vl_logic_vector(31 downto 0);
        oFREE_SET_IRQ_MODE: out    vl_logic;
        oFREE_CLR_IRQ_MODE: out    vl_logic;
        oFREE_CACHE_FLUSH: out    vl_logic;
        oFREE_TLB_FLUSH : out    vl_logic;
        iINTERRUPT_LOCK : in     vl_logic;
        iINTERRUPT_LDST_LOCK: in     vl_logic;
        iSYSREG_SPR     : in     vl_logic_vector(31 downto 0);
        iSYSREG_TIDR    : in     vl_logic_vector(31 downto 0);
        iSYSREG_TISR    : in     vl_logic_vector(31 downto 0);
        iSYSREG_PSR     : in     vl_logic_vector(31 downto 0);
        iSYSREG_PPSR    : in     vl_logic_vector(31 downto 0);
        iSYSREG_PCR     : in     vl_logic_vector(31 downto 0);
        iSYSREG_PPCR    : in     vl_logic_vector(31 downto 0);
        iSYSREG_IDTR    : in     vl_logic_vector(31 downto 0);
        oSYSREG_SPR_WRITE: out    vl_logic;
        oSYSREG_SPR     : out    vl_logic_vector(31 downto 0);
        oLDST_USE       : out    vl_logic;
        oLDST_REQ       : out    vl_logic;
        iLDST_BUSY      : in     vl_logic;
        oLDST_ORDER     : out    vl_logic_vector(1 downto 0);
        oLDST_RW        : out    vl_logic;
        oLDST_TID       : out    vl_logic_vector(13 downto 0);
        oLDST_MMUMOD    : out    vl_logic_vector(1 downto 0);
        oLDST_PDT       : out    vl_logic_vector(31 downto 0);
        oLDST_ADDR      : out    vl_logic_vector(31 downto 0);
        oLDST_DATA      : out    vl_logic_vector(31 downto 0);
        iLDST_REQ       : in     vl_logic;
        iLDST_DATA      : in     vl_logic_vector(31 downto 0);
        oIO_IRQ_CONFIG_TABLE_REQ: out    vl_logic;
        oIO_IRQ_CONFIG_TABLE_ENTRY: out    vl_logic_vector(5 downto 0);
        oIO_IRQ_CONFIG_TABLE_FLAG_MASK: out    vl_logic;
        oIO_IRQ_CONFIG_TABLE_FLAG_VALID: out    vl_logic;
        oIO_IRQ_CONFIG_TABLE_FLAG_LEVEL: out    vl_logic_vector(1 downto 0);
        oICT_REQ        : out    vl_logic;
        oICT_ENTRY      : out    vl_logic_vector(5 downto 0);
        oICT_CONF_MASK  : out    vl_logic;
        oICT_CONF_VALID : out    vl_logic;
        oICT_CONF_LEVEL : out    vl_logic_vector(1 downto 0);
        iEXCEPT_JUMP    : in     vl_logic;
        iEXCEPT_JUMP_ADDR: in     vl_logic_vector(31 downto 0);
        iEXCEPT_IDTS    : in     vl_logic;
        iEXCEPT_IDTS_ADDR: in     vl_logic_vector(31 downto 0);
        iEXCEPT_IB      : in     vl_logic;
        iEXCEPT_IB_ADDR : in     vl_logic_vector(31 downto 0);
        iEXCEPT_PDTS    : in     vl_logic;
        iEXCEPT_IRQ_REQ : in     vl_logic;
        iEXCEPT_IRQ_NUM : in     vl_logic_vector(6 downto 0);
        iEXCEPT_IRQ_FI0R: in     vl_logic_vector(31 downto 0);
        oEXCEPT_IRQ_ACK : out    vl_logic;
        oEXCEPT_IRQ_BUSY: out    vl_logic
    );
end exception_manager;
