library verilog;
use verilog.vl_types.all;
entity memory_pipe_arbiter is
    port(
        iCLOCK          : in     vl_logic;
        inRESET         : in     vl_logic;
        iDATA_REQ       : in     vl_logic;
        oDATA_LOCK      : out    vl_logic;
        iDATA_ORDER     : in     vl_logic_vector(1 downto 0);
        iDATA_MASK      : in     vl_logic_vector(3 downto 0);
        iDATA_RW        : in     vl_logic;
        iDATA_TID       : in     vl_logic_vector(13 downto 0);
        iDATA_MMUMOD    : in     vl_logic_vector(1 downto 0);
        iDATA_MMUPS     : in     vl_logic_vector(2 downto 0);
        iDATA_PDT       : in     vl_logic_vector(31 downto 0);
        iDATA_ADDR      : in     vl_logic_vector(31 downto 0);
        iDATA_DATA      : in     vl_logic_vector(31 downto 0);
        oDATA_REQ       : out    vl_logic;
        iDATA_BUSY      : in     vl_logic;
        oDATA_DATA      : out    vl_logic_vector(63 downto 0);
        oDATA_MMU_FLAGS : out    vl_logic_vector(23 downto 0);
        iINST_REQ       : in     vl_logic;
        oINST_LOCK      : out    vl_logic;
        iINST_MMUMOD    : in     vl_logic_vector(1 downto 0);
        iINST_MMUPS     : in     vl_logic_vector(2 downto 0);
        iINST_PDT       : in     vl_logic_vector(31 downto 0);
        iINST_ADDR      : in     vl_logic_vector(31 downto 0);
        oINST_REQ       : out    vl_logic;
        iINST_BUSY      : in     vl_logic;
        oINST_DATA      : out    vl_logic_vector(63 downto 0);
        oINST_MMU_FLAGS : out    vl_logic_vector(23 downto 0);
        oMEMORY_REQ     : out    vl_logic;
        iMEMORY_LOCK    : in     vl_logic;
        oMEMORY_DATA_STORE_ACK: out    vl_logic;
        oMEMORY_MMU_MODE: out    vl_logic_vector(1 downto 0);
        oMEMORY_MMU_PS  : out    vl_logic_vector(2 downto 0);
        oMEMORY_PDT     : out    vl_logic_vector(31 downto 0);
        oMEMORY_ORDER   : out    vl_logic_vector(1 downto 0);
        oMEMORY_MASK    : out    vl_logic_vector(3 downto 0);
        oMEMORY_RW      : out    vl_logic;
        oMEMORY_ADDR    : out    vl_logic_vector(31 downto 0);
        oMEMORY_DATA    : out    vl_logic_vector(31 downto 0);
        iMEMORY_VALID   : in     vl_logic;
        oMEMORY_BUSY    : out    vl_logic;
        iMEMORY_STORE_ACK: in     vl_logic;
        iMEMORY_DATA    : in     vl_logic_vector(63 downto 0);
        iMEMORY_MMU_FLAGS: in     vl_logic_vector(23 downto 0)
    );
end memory_pipe_arbiter;
