library verilog;
use verilog.vl_types.all;
entity dispatch is
    generic(
        CORE_ID         : integer := 0
    );
    port(
        iCLOCK          : in     vl_logic;
        inRESET         : in     vl_logic;
        iFREE_REGISTER_LOCK: in     vl_logic;
        iFREE_PIPELINE_STOP: in     vl_logic;
        iFREE_REFRESH   : in     vl_logic;
        oEXCEPTION_LOCK : out    vl_logic;
        iSYSREGINFO_IOSR_VALID: in     vl_logic;
        iSYSREGINFO_IOSR: in     vl_logic_vector(31 downto 0);
        iFREE_SYSREG_SET_IRQ_MODE: in     vl_logic;
        iFREE_SYSREG_CLR_IRQ_MODE: in     vl_logic;
        iFREE_PPCR_SET  : in     vl_logic;
        iFREE_PPCR      : in     vl_logic_vector(31 downto 0);
        iFREE_FI0R_SET  : in     vl_logic;
        iFREE_FI0R      : in     vl_logic_vector(31 downto 0);
        iSYSREG_FLAGR   : in     vl_logic_vector(31 downto 0);
        oSYSREG_PCR     : out    vl_logic_vector(31 downto 0);
        oSYSREG_IDTR    : out    vl_logic_vector(31 downto 0);
        oSYSREG_TISR    : out    vl_logic_vector(31 downto 0);
        oSYSREG_TIDR    : out    vl_logic_vector(31 downto 0);
        oSYSREG_PSR     : out    vl_logic_vector(31 downto 0);
        oSYSREG_PPSR    : out    vl_logic_vector(31 downto 0);
        oSYSREG_PPCR    : out    vl_logic_vector(31 downto 0);
        oSYSREG_SPR     : out    vl_logic_vector(31 downto 0);
        iPREVIOUS_VALID : in     vl_logic;
        iPREVIOUS_FAULT_PAGEFAULT: in     vl_logic;
        iPREVIOUS_FAULT_PRIVILEGE_ERROR: in     vl_logic;
        iPREVIOUS_FAULT_INVALID_INST: in     vl_logic;
        iPREVIOUS_PAGING_ENA: in     vl_logic;
        iPREVIOUS_KERNEL_ACCESS: in     vl_logic;
        iPREVIOUS_BRANCH_PREDICT: in     vl_logic;
        iPREVIOUS_BRANCH_PREDICT_ADDR: in     vl_logic_vector(31 downto 0);
        iPREVIOUS_SOURCE0_ACTIVE: in     vl_logic;
        iPREVIOUS_SOURCE1_ACTIVE: in     vl_logic;
        iPREVIOUS_SOURCE0_SYSREG: in     vl_logic;
        iPREVIOUS_SOURCE1_SYSREG: in     vl_logic;
        iPREVIOUS_ADV_ACTIVE: in     vl_logic;
        iPREVIOUS_DESTINATION_SYSREG: in     vl_logic;
        iPREVIOUS_DESTINATION: in     vl_logic_vector(4 downto 0);
        iPREVIOUS_WRITEBACK: in     vl_logic;
        iPREVIOUS_FLAGS_WRITEBACK: in     vl_logic;
        iPREVIOUS_CMD   : in     vl_logic_vector(4 downto 0);
        iPREVIOUS_CC_AFE: in     vl_logic_vector(3 downto 0);
        iPREVIOUS_SOURCE0: in     vl_logic_vector(4 downto 0);
        iPREVIOUS_SOURCE1: in     vl_logic_vector(31 downto 0);
        iPREVIOUS_ADV_DATA: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_SOURCE0_FLAGS: in     vl_logic;
        iPREVIOUS_SOURCE1_IMM: in     vl_logic;
        iPREVIOUS_EX_SYS_REG: in     vl_logic;
        iPREVIOUS_EX_SYS_LDST: in     vl_logic;
        iPREVIOUS_EX_LOGIC: in     vl_logic;
        iPREVIOUS_EX_SHIFT: in     vl_logic;
        iPREVIOUS_EX_ADDER: in     vl_logic;
        iPREVIOUS_EX_MUL: in     vl_logic;
        iPREVIOUS_EX_SDIV: in     vl_logic;
        iPREVIOUS_EX_UDIV: in     vl_logic;
        iPREVIOUS_EX_LDST: in     vl_logic;
        iPREVIOUS_EX_BRANCH: in     vl_logic;
        iPREVIOUS_PC    : in     vl_logic_vector(31 downto 0);
        oPREVIOUS_LOCK  : out    vl_logic;
        oNEXT_VALID     : out    vl_logic;
        oNEXT_FAULT_PAGEFAULT: out    vl_logic;
        oNEXT_FAULT_PRIVILEGE_ERROR: out    vl_logic;
        oNEXT_FAULT_INVALID_INST: out    vl_logic;
        oNEXT_PAGING_ENA: out    vl_logic;
        oNEXT_KERNEL_ACCESS: out    vl_logic;
        oNEXT_BRANCH_PREDICT: out    vl_logic;
        oNEXT_BRANCH_PREDICT_ADDR: out    vl_logic_vector(31 downto 0);
        oNEXT_SYSREG_PSR: out    vl_logic_vector(31 downto 0);
        oNEXT_SYSREG_TIDR: out    vl_logic_vector(31 downto 0);
        oNEXT_SYSREG_PDTR: out    vl_logic_vector(31 downto 0);
        oNEXT_DESTINATION_SYSREG: out    vl_logic;
        oNEXT_DESTINATION: out    vl_logic_vector(4 downto 0);
        oNEXT_WRITEBACK : out    vl_logic;
        oNEXT_FLAGS_WRITEBACK: out    vl_logic;
        oNEXT_CMD       : out    vl_logic_vector(4 downto 0);
        oNEXT_CC_AFE    : out    vl_logic_vector(3 downto 0);
        oNEXT_SPR       : out    vl_logic_vector(31 downto 0);
        oNEXT_SOURCE0   : out    vl_logic_vector(31 downto 0);
        oNEXT_SOURCE1   : out    vl_logic_vector(31 downto 0);
        oNEXT_ADV_DATA  : out    vl_logic_vector(5 downto 0);
        oNEXT_SOURCE0_POINTER: out    vl_logic_vector(4 downto 0);
        oNEXT_SOURCE1_POINTER: out    vl_logic_vector(4 downto 0);
        oNEXT_SOURCE0_SYSREG: out    vl_logic;
        oNEXT_SOURCE1_SYSREG: out    vl_logic;
        oNEXT_SOURCE1_IMM: out    vl_logic;
        oNEXT_SOURCE0_FLAGS: out    vl_logic;
        oNEXT_ADV_ACTIVE: out    vl_logic;
        oNEXT_EX_SYS_REG: out    vl_logic;
        oNEXT_EX_SYS_LDST: out    vl_logic;
        oNEXT_EX_LOGIC  : out    vl_logic;
        oNEXT_EX_SHIFT  : out    vl_logic;
        oNEXT_EX_ADDER  : out    vl_logic;
        oNEXT_EX_MUL    : out    vl_logic;
        oNEXT_EX_SDIV   : out    vl_logic;
        oNEXT_EX_UDIV   : out    vl_logic;
        oNEXT_EX_LDST   : out    vl_logic;
        oNEXT_EX_BRANCH : out    vl_logic;
        oNEXT_PC        : out    vl_logic_vector(31 downto 0);
        iNEXT_LOCK      : in     vl_logic;
        iWB_VALID       : in     vl_logic;
        iWB_DATA        : in     vl_logic_vector(31 downto 0);
        iWB_DESTINATION : in     vl_logic_vector(4 downto 0);
        iWB_DESTINATION_SYSREG: in     vl_logic;
        iWB_WRITEBACK   : in     vl_logic;
        iWB_SPR_WRITEBACK: in     vl_logic;
        iWB_SPR         : in     vl_logic_vector(31 downto 0);
        iWB_PC          : in     vl_logic_vector(31 downto 0);
        iWB_BRANCH      : in     vl_logic;
        iWB_BRANCH_PC   : in     vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR0: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR1: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR2: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR3: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR4: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR5: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR6: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR7: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR8: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR9: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR10: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR11: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR12: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR13: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR14: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR15: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR16: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR17: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR18: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR19: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR20: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR21: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR22: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR23: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR24: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR25: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR26: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR27: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR28: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR29: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR30: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_GR31: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_SPR: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_PCR: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_PPCR: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_PSR: out    vl_logic_vector(31 downto 0);
        oDEBUG_REG_OUT_PPSR: out    vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CORE_ID : constant is 1;
end dispatch;
