library verilog;
use verilog.vl_types.all;
entity mist1032isa is
    port(
        iCORE_CLOCK     : in     vl_logic;
        iBUS_CLOCK      : in     vl_logic;
        iDPS_CLOCK      : in     vl_logic;
        inRESET         : in     vl_logic;
        oSCI_TXD        : out    vl_logic;
        iSCI_RXD        : in     vl_logic;
        oMEMORY_REQ     : out    vl_logic;
        iMEMORY_LOCK    : in     vl_logic;
        oMEMORY_ORDER   : out    vl_logic_vector(1 downto 0);
        oMEMORY_MASK    : out    vl_logic_vector(3 downto 0);
        oMEMORY_RW      : out    vl_logic;
        oMEMORY_ADDR    : out    vl_logic_vector(31 downto 0);
        oMEMORY_DATA    : out    vl_logic_vector(31 downto 0);
        iMEMORY_VALID   : in     vl_logic;
        oMEMORY_BUSY    : out    vl_logic;
        iMEMORY_DATA    : in     vl_logic_vector(63 downto 0);
        oGCI_REQ        : out    vl_logic;
        iGCI_BUSY       : in     vl_logic;
        oGCI_RW         : out    vl_logic;
        oGCI_ADDR       : out    vl_logic_vector(31 downto 0);
        oGCI_DATA       : out    vl_logic_vector(31 downto 0);
        iGCI_REQ        : in     vl_logic;
        oGCI_BUSY       : out    vl_logic;
        iGCI_DATA       : in     vl_logic_vector(31 downto 0);
        iGCI_IRQ_REQ    : in     vl_logic;
        iGCI_IRQ_NUM    : in     vl_logic_vector(5 downto 0);
        oGCI_IRQ_ACK    : out    vl_logic;
        oIO_IRQ_CONFIG_TABLE_REQ: out    vl_logic;
        oIO_IRQ_CONFIG_TABLE_ENTRY: out    vl_logic_vector(5 downto 0);
        oIO_IRQ_CONFIG_TABLE_FLAG_MASK: out    vl_logic;
        oIO_IRQ_CONFIG_TABLE_FLAG_VALID: out    vl_logic;
        oIO_IRQ_CONFIG_TABLE_FLAG_LEVEL: out    vl_logic_vector(1 downto 0);
        oDEBUG_PC       : out    vl_logic_vector(31 downto 0);
        oDEBUG0         : out    vl_logic_vector(31 downto 0);
        iDEBUG_UART_RXD : in     vl_logic;
        oDEBUG_UART_TXD : out    vl_logic;
        iDEBUG_PARA_REQ : in     vl_logic;
        oDEBUG_PARA_BUSY: out    vl_logic;
        iDEBUG_PARA_CMD : in     vl_logic_vector(7 downto 0);
        iDEBUG_PARA_DATA: in     vl_logic_vector(31 downto 0);
        oDEBUG_PARA_VALID: out    vl_logic;
        iDEBUG_PARA_BUSY: in     vl_logic;
        oDEBUG_PARA_ERROR: out    vl_logic;
        oDEBUG_PARA_DATA: out    vl_logic_vector(31 downto 0)
    );
end mist1032isa;
