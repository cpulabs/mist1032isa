library verilog;
use verilog.vl_types.all;
entity load_store_pipe_arbiter is
    port(
        oLDST_REQ       : out    vl_logic;
        iLDST_BUSY      : in     vl_logic;
        oLDST_ORDER     : out    vl_logic_vector(1 downto 0);
        oLDST_MASK      : out    vl_logic_vector(3 downto 0);
        oLDST_RW        : out    vl_logic;
        oLDST_TID       : out    vl_logic_vector(13 downto 0);
        oLDST_MMUMOD    : out    vl_logic_vector(1 downto 0);
        oLDST_MMUPS     : out    vl_logic_vector(2 downto 0);
        oLDST_PDT       : out    vl_logic_vector(31 downto 0);
        oLDST_ADDR      : out    vl_logic_vector(31 downto 0);
        oLDST_DATA      : out    vl_logic_vector(31 downto 0);
        iLDST_VALID     : in     vl_logic;
        iLDST_MMU_FLAGS : in     vl_logic_vector(11 downto 0);
        iLDST_DATA      : in     vl_logic_vector(31 downto 0);
        iUSE_SEL        : in     vl_logic;
        iEXE_REQ        : in     vl_logic;
        oEXE_BUSY       : out    vl_logic;
        iEXE_ORDER      : in     vl_logic_vector(1 downto 0);
        iEXE_MASK       : in     vl_logic_vector(3 downto 0);
        iEXE_RW         : in     vl_logic;
        iEXE_TID        : in     vl_logic_vector(13 downto 0);
        iEXE_MMUMOD     : in     vl_logic_vector(1 downto 0);
        iEXE_MMUPS      : in     vl_logic_vector(2 downto 0);
        iEXE_PDT        : in     vl_logic_vector(31 downto 0);
        iEXE_ADDR       : in     vl_logic_vector(31 downto 0);
        iEXE_DATA       : in     vl_logic_vector(31 downto 0);
        oEXE_REQ        : out    vl_logic;
        oEXE_MMU_FLAGS  : out    vl_logic_vector(11 downto 0);
        oEXE_DATA       : out    vl_logic_vector(31 downto 0);
        iEXCEPT_REQ     : in     vl_logic;
        oEXCEPT_BUSY    : out    vl_logic;
        iEXCEPT_ORDER   : in     vl_logic_vector(1 downto 0);
        iEXCEPT_RW      : in     vl_logic;
        iEXCEPT_TID     : in     vl_logic_vector(13 downto 0);
        iEXCEPT_MMUMOD  : in     vl_logic_vector(1 downto 0);
        iEXCEPT_MMUPS   : in     vl_logic_vector(2 downto 0);
        iEXCEPT_PDT     : in     vl_logic_vector(31 downto 0);
        iEXCEPT_ADDR    : in     vl_logic_vector(31 downto 0);
        iEXCEPT_DATA    : in     vl_logic_vector(31 downto 0);
        oEXCEPT_REQ     : out    vl_logic;
        oEXCEPT_DATA    : out    vl_logic_vector(31 downto 0)
    );
end load_store_pipe_arbiter;
